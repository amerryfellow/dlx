package alu_types is
	type TYPE_OP is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, LSL, LSR, LRL, LRR);
end types;
