package CONSTANTS is
   constant INVERTER_DELAY : time := 0.1 ns;
   constant NAND1_DELAY : time := 0.2 ns;
   constant NDDELAYRISE : time := 0.6 ns;
   constant NDDELAYFALL : time := 0.4 ns;
   constant NOR_DELAY : time := 0.2 ns;
   constant RIPPLECARRYADDER_DELAY_S : time := 1 ns;
   constant DIPPLECARRYADDER_DELAY_C : time := 2 ns;
   constant NumBit : integer := 4;	
   constant TP_MUX : time := 0.5 ns; 	
end CONSTANTS;
