library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;
use WORK.alu_types.all;

-- Behavioral

entity SUMGENERATOR is
	generic(
		NBIT:	integer	:= NSUMG; --32,64 
		NCSB:	integer	:= NCSUMG --8,16
	);
	port (
		A:	in	std_logic_vector(NBIT-1 downto 0);
		B:	in	std_logic_vector(NBIT-1 downto 0);
		Ci:	in	std_logic_vector(NCSB-1 downto 0);
		S:	out	std_logic_vector(NBIT-1 downto 0)
	);
end SUMGENERATOR;

-- Architectures

architecture structural of SUMGENERATOR is
	component CSB 
		generic(
			N:	integer	:= NCSBLOCK -- 4
		);
		port (
			A:	in	std_logic_vector(N-1 downto 0);
			B:	in	std_logic_vector(N-1 downto 0);
			Ci:	in	std_logic;
			S:	out	std_logic_vector(N-1 downto 0)
		);
	end component;
	
begin
	-- For NCSBLOCK and others constants refer to P4ADDER_constants file.
	-- This structural architecture generates (NCSB - 1) carry selects block of NCSBLOCK bits,
	-- which is the number of carry bits generated by the sparse tree, plus 1, that is the carry in.

	CS: for i in 0 to NCSB-1 generate
		CSBX: CSB
			port map(
				A(((i*NCSBLOCK)+NCSBLOCK-1) downto i*NCSBLOCK),
				B(((i*NCSBLOCK)+NCSBLOCK-1) downto i*NCSBLOCK),
				Ci(i),
				S(((i*NCSBLOCK)+NCSBLOCK-1) downto i*NCSBLOCK)
			);
	end generate;
end structural;

