ripplecarryadder/rca_generic.vhd