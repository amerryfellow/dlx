package GENERICS is
   constant NumBit : integer := 8;		
end GENERICS;
