package CONSTANTS is
   constant IVDELAY : time := 0.1 ns;
   constant NDDELAY : time := 0.2 ns;
   constant NDDELAYRISE : time := 0.6 ns;
   constant NDDELAYFALL : time := 0.4 ns;
   constant NRDELAY : time := 0.2 ns;
   constant DRCAS : time := 1 ps;
   constant DRCAC : time := 2 ps;
   constant DFAS: time := 0.5 ps;
   constant DFAC: time := 1 ps;
   constant NumBit : integer := 64;	
   constant TP_MUX : time := 0.5 ps; 	
end CONSTANTS;
