mux/mux.vhd