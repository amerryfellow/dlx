package CONSTANTS is
   constant adderBits : integer := 64;
   constant multiplierBits : integer := 8;
   constant defaultBits : integer := 8;
   constant TP_MUX : time := 0.5 ps;
end CONSTANTS;
